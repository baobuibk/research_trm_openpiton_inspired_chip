// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// Author: Michael Schaffner <schaffner@iis.ee.ethz.ch>, ETH Zurich
// Date: 19.03.2017
// Description: Ariane Top-level wrapper to break out SV structs to logic vectors.

`define NrMaxRules_V 16
module ariane_verilog_wrap #(
  parameter int unsigned CORE_ADDR                           = 1,
  parameter int unsigned               RASDepth              = 2,
  parameter int unsigned               BTBEntries            = 32,
  parameter int unsigned               BHTEntries            = 128,
  // debug module base address
  parameter logic [63:0]               DmBaseAddress         = 64'h0,
  // swap endianess in l15 adapter
  parameter bit                        SwapEndianess         = 1,
  // PMA configuration
  // idempotent region
  parameter int unsigned               NrNonIdempotentRules  =  0,
  parameter logic [`NrMaxRules_V*64-1:0]  NonIdempotentAddrBase = '0,
  parameter logic [`NrMaxRules_V*64-1:0]  NonIdempotentLength   = '0,
  // executable regions
  parameter int unsigned               NrExecuteRegionRules  =  0,
  parameter logic [`NrMaxRules_V*64-1:0]  ExecuteRegionAddrBase = '0,
  parameter logic [`NrMaxRules_V*64-1:0]  ExecuteRegionLength   = '0,
  // cacheable regions
  parameter int unsigned               NrCachedRegionRules   =  0,
  parameter logic [`NrMaxRules_V*64-1:0]  CachedRegionAddrBase  = '0,
  parameter logic [`NrMaxRules_V*64-1:0]  CachedRegionLength    = '0
) (
  input                       clk_i,
  input                       reset_l,      // this is an openpiton-specific name, do not change (hier. paths in TB use this)
  output                      spc_grst_l,   // this is an openpiton-specific name, do not change (hier. paths in TB use this)
  // Core ID, Cluster ID and boot address are considered more or less static
  input  [63:0]               boot_addr_i,  // reset boot address
  input  [63:0]               hart_id_i,    // hart id in a multicore environment (reflected in a CSR)
  // Interrupt inputs
  input  [1:0]                irq_i,        // level sensitive IR lines, mip & sip (async)
  input                       ipi_i,        // inter-processor interrupts (async)
  // Timer facilities
  input                       time_irq_i,   // timer interrupt in (async)
  input                       debug_req_i,  // debug request (async)

`ifdef PITON_ARIANE
  // L15 (memory side)
  output [$size(wt_cache_pkg::l15_req_t)-1:0]  l15_req_o,
  input  [$size(wt_cache_pkg::l15_rtrn_t)-1:0] l15_rtrn_i
`else
  // AXI (memory side)
  output [$size(ariane_axi::req_t)-1:0]             axi_req_o,
  input  [$size(ariane_axi::resp_t)-1:0]            axi_resp_i
`endif
 );

// assign bitvector to packed struct and vice versa
`ifdef PITON_ARIANE
  // L15 (memory side)
  wt_cache_pkg::l15_req_t  l15_req;
  wt_cache_pkg::l15_rtrn_t l15_rtrn;

  assign l15_req_o = l15_req;
  assign l15_rtrn  = l15_rtrn_i;
`else
  ariane_axi::req_t             axi_req;
  ariane_axi::resp_t            axi_resp;

  assign axi_req_o = axi_req;
  assign axi_resp  = axi_resp_i;
`endif


  /////////////////////////////
  // Core wakeup mechanism
  /////////////////////////////

  logic [15:0] wake_up_cnt_d, wake_up_cnt_q;
  logic rst_n;

  assign wake_up_cnt_d = (wake_up_cnt_q[$high(wake_up_cnt_q)]) ? wake_up_cnt_q : wake_up_cnt_q + 1;

  always_ff @(posedge clk_i or negedge reset_l) begin : p_regs
    if(~reset_l) begin
      wake_up_cnt_q <= 0;
    end else begin
      wake_up_cnt_q <= wake_up_cnt_d;
    end
  end

  // reset gate this
  //assign rst_n = wake_up_cnt_q[$high(wake_up_cnt_q)] & reset_l;
  assign rst_n = wake_up_cnt_q > 5018 ? 1 : 0;

  /////////////////////////////
  // synchronizers
  /////////////////////////////

  logic [1:0] irq;
  logic ipi, time_irq, debug_req;

  // reset synchronization
  synchronizer i_sync (
    .clk         ( clk_i      ),
    .presyncdata ( rst_n      ),
    .syncdata    ( spc_grst_l )
  );

  // interrupts
  for (genvar k=0; k<$size(irq_i); k++) begin
    synchronizer i_irq_sync (
      .clk         ( clk_i      ),
      .presyncdata ( irq_i[k]   ),
      .syncdata    ( irq[k]     )
    );
  end

  synchronizer i_ipi_sync (
    .clk         ( clk_i      ),
    .presyncdata ( ipi_i      ),
    .syncdata    ( ipi        )
  );

  synchronizer i_timer_sync (
    .clk         ( clk_i      ),
    .presyncdata ( time_irq_i ),
    .syncdata    ( time_irq   )
  );

  synchronizer i_debug_sync (
    .clk         ( clk_i       ),
    .presyncdata ( debug_req_i ),
    .syncdata    ( debug_req   )
  );

  /////////////////////////////
  // ariane instance
  /////////////////////////////

  localparam ariane_pkg::ariane_cfg_t ArianeOpenPitonCfg = '{
    RASDepth:              RASDepth,
    BTBEntries:            BTBEntries,
    BHTEntries:            BHTEntries,
    // idempotent region
    NrNonIdempotentRules:  NrNonIdempotentRules,
    NonIdempotentAddrBase: NonIdempotentAddrBase,
    NonIdempotentLength:   NonIdempotentLength,
    NrExecuteRegionRules:  NrExecuteRegionRules,
    ExecuteRegionAddrBase: ExecuteRegionAddrBase,
    ExecuteRegionLength:   ExecuteRegionLength,
    // cached region
    NrCachedRegionRules:   NrCachedRegionRules,
    CachedRegionAddrBase:  CachedRegionAddrBase,
    CachedRegionLength:    CachedRegionLength,
    // cache config
    Axi64BitCompliant:     1'b0,
    SwapEndianess:         SwapEndianess,
    // debug
    DmBaseAddress:         DmBaseAddress
  };

  ariane #(
    .CORE_ADDR(CORE_ADDR),
    .ArianeCfg ( ArianeOpenPitonCfg )
  ) ariane (
    .clk_i       ( clk_i      ),
    .rst_ni      ( spc_grst_l ),
    .boot_addr_i              ,// constant
    .hart_id_i                ,// constant
    .irq_i       ( irq        ),
    .ipi_i       ( ipi        ),
    .time_irq_i  ( time_irq   ),
    .debug_req_i ( debug_req  ),
`ifdef PITON_ARIANE
    .l15_req_o   ( l15_req   ),
    .l15_rtrn_i  ( l15_rtrn  )
`else
    .axi_req_o   ( axi_req   ),
    .axi_resp_i  ( axi_resp  )
`endif
  );

endmodule // ariane_verilog_wrap
